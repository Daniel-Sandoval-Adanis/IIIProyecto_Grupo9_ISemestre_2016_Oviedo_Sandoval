`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:05:23 05/30/2016 
// Design Name: 
// Module Name:    Controlador_VGA 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Controlador_VGA(
	 input wire [7:0] dato2,dato0, 
	 input wire crontermino,
	 input wire [3:0] dig0, dig1,dig2, dig3,dig4, dig5,dig6, dig7,dig8, dig9,dig10, dig11,dig12, dig13,dig14, dig15,dig16, dig17,
	 input wire clk,reset,
	 output wire hsync, vsync,
    output wire [7:0] text_rgb
    );


endmodule
